
/********************************************************
** Waveform Generator and Radar Control Blocks: 64-127
********************************************************/
localparam [7:0] SR_CH_COUNTER_ADDR = 64;
localparam [7:0] SR_CH_TUNING_COEF_ADDR = 65;
localparam [7:0] SR_CH_FREQ_OFFSET_ADDR = 66;
localparam [7:0] SR_AWG_CTRL_WORD_ADDR = 67;

localparam [7:0] SR_PRF_INT_ADDR = 68;
localparam [7:0] SR_PRF_FRAC_ADDR = 69;
localparam [7:0] SR_ADC_SAMPLE_ADDR = 70;
